module spitb ;
  
  reg clk1;
  reg sclk1;
  wire dout1;
  reg din1;
  wire [4:0] count1;
  wire cs1;
  wire [1:0] rst1;
  
  
  initial begin 
    
    $dumpfile("dump.vcd");
    $dumpvars(1);
    
    clk1<=0;#10; 
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=0;#10; 
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=0;#10; 
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
    clk1<=1;#10;
    clk1<=0;#10;
  end
  
  spi inter(.clk(clk1), .sclk(sclk1), .din(din1), .dout(dout1), .cs(cs1), .count(count1), .rst(rst1));
  
    
endmodule